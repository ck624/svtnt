/****************************************************************************
 * svtnt_pkg.sv
 ****************************************************************************/

/**
 * Package: svtnt_pkg
 * 
 * TODO: Add package documentation
 */
package svtnt_pkg;

	import "SVTNT" __svtnt_display=function void \$display (string fmt, ...);


endpackage


